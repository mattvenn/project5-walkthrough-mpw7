VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO rgb_mixer
  CLASS BLOCK ;
  FOREIGN rgb_mixer ;
  ORIGIN 0.000 0.000 ;
  SIZE 250.000 BY 250.000 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 122.440 250.000 123.040 ;
    END
  END clk
  PIN enc0_a
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.310 246.000 3.590 250.000 ;
    END
  END enc0_a
  PIN enc0_b
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 187.040 250.000 187.640 ;
    END
  END enc0_b
  PIN enc1_a
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.810 0.000 245.090 4.000 ;
    END
  END enc1_a
  PIN enc1_b
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.670 246.000 125.950 250.000 ;
    END
  END enc1_b
  PIN enc2_a
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END enc2_a
  PIN enc2_b
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.630 0.000 183.910 4.000 ;
    END
  END enc2_b
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.270 0.000 61.550 4.000 ;
    END
  END io_oeb[0]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.850 246.000 187.130 250.000 ;
    END
  END io_oeb[1]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.240 4.000 61.840 ;
    END
  END io_oeb[2]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 125.840 4.000 126.440 ;
    END
  END io_oeb[3]
  PIN pwm0_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.030 246.000 248.310 250.000 ;
    END
  END pwm0_out
  PIN pwm1_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.450 0.000 122.730 4.000 ;
    END
  END pwm1_out
  PIN pwm2_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 190.440 4.000 191.040 ;
    END
  END pwm2_out
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.490 246.000 64.770 250.000 ;
    END
  END reset
  PIN sync
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 57.840 250.000 58.440 ;
    END
  END sync
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 236.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 236.880 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 236.880 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 244.260 236.725 ;
      LAYER met1 ;
        RECT 0.070 10.640 248.330 236.880 ;
      LAYER met2 ;
        RECT 0.100 245.720 3.030 246.570 ;
        RECT 3.870 245.720 64.210 246.570 ;
        RECT 65.050 245.720 125.390 246.570 ;
        RECT 126.230 245.720 186.570 246.570 ;
        RECT 187.410 245.720 247.750 246.570 ;
        RECT 0.100 4.280 248.300 245.720 ;
        RECT 0.650 4.000 60.990 4.280 ;
        RECT 61.830 4.000 122.170 4.280 ;
        RECT 123.010 4.000 183.350 4.280 ;
        RECT 184.190 4.000 244.530 4.280 ;
        RECT 245.370 4.000 248.300 4.280 ;
      LAYER met3 ;
        RECT 4.000 191.440 246.000 236.805 ;
        RECT 4.400 190.040 246.000 191.440 ;
        RECT 4.000 188.040 246.000 190.040 ;
        RECT 4.000 186.640 245.600 188.040 ;
        RECT 4.000 126.840 246.000 186.640 ;
        RECT 4.400 125.440 246.000 126.840 ;
        RECT 4.000 123.440 246.000 125.440 ;
        RECT 4.000 122.040 245.600 123.440 ;
        RECT 4.000 62.240 246.000 122.040 ;
        RECT 4.400 60.840 246.000 62.240 ;
        RECT 4.000 58.840 246.000 60.840 ;
        RECT 4.000 57.440 245.600 58.840 ;
        RECT 4.000 10.715 246.000 57.440 ;
  END
END rgb_mixer
END LIBRARY

